module main

import server

fn main() {
    server.run()
}

