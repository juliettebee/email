module main

import smtp_server 

fn main() {
    smtp_server.start()
}

